module ALU_Deco(
    input logic [6:0]   op,
    input logic [2:0]   funct3,
    input logic         funct7_5,
    input logic [1:0]   ALUOp

    output logic [2:0]  ALUControl
)

always_comb
    case (ALUOp)
        2'b00: ALUControl = 3'b000;
        2'b01: ALUControl = 3'b001;
        2'b10: 
            case(funct3)
                3'b000: 
                    if op[5] & funct7_5 == 1'b1
                        ALUControl = 3'b001;
                    else
                        ALUControl = 3'b000;
        
                3'b010: ALUControl = 3'b101;
                3'b110: ALUControl = 3'b011;
                3'b111: ALUControl = 3'b010;
                default: ALUControl = 3'b000;
            endcase
        default: ALUControl = 3'b000;
    endcase
        
endmodule